`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NUS
// Engineer: Shahzor Ahmad, Rajesh C Panicker
// 
// Create Date: 27.09.2016 10:59:44
// Design Name: 
// Module Name: MCycle
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
/* 
----------------------------------------------------------------------------------
--	(c) Shahzor Ahmad, Rajesh C Panicker
--	License terms :
--	You are free to use this code as long as you
--		(i) DO NOT post it on any public repository;
--		(ii) use it only for educational purposes;
--		(iii) accept the responsibility to ensure that your implementation does not violate any intellectual property of ARM Holdings or other entities.
--		(iv) accept that the program is provided "as is" without warranty of any kind or assurance regarding its suitability for any particular purpose;
--		(v) send an email to rajesh.panicker@ieee.org briefly mentioning its use (except when used for the course CG3207 at the National University of Singapore);
--		(vi) retain this notice in this file or any files derived from this.
----------------------------------------------------------------------------------
*/

module MCycle

    #(parameter width = 4) // Keep this at 4 to verify your algorithms with 4 bit numbers (easier). When using MCycle as a component in ARM, generic map it to 32.
    (
        input CLK,
        input RESET, // Connect this to the reset of the ARM processor.
        input Start, // Multi-cycle Enable. The control unit should assert this when an instruction with a multi-cycle operation is detected.
        input [1:0] MCycleOp, // Multi-cycle Operation. "00" for signed multiplication, "01" for unsigned multiplication, "10" for signed division, "11" for unsigned division. Generated by Control unit
        input [width-1:0] Operand1, // Multiplicand / Dividend
        input [width-1:0] Operand2, // Multiplier / Divisor
        output reg [width-1:0] Result1, // LSW of Product / Quotient
        output reg [width-1:0] Result2, // MSW of Product / Remainder
        output reg Busy // Set immediately when Start is set. Cleared when the Results become ready. This bit can be used to stall the processor while multi-cycle operations are on.
    );
    
// use the Busy signal to reset WE_PC to 0 in ARM.v (aka "freeze" PC). The two signals are complements of each other
// since the IDLE_PROCESS is combinational, instantaneously asserts Busy once Start is asserted
  
    parameter IDLE = 1'b0 ;  // will cause a warning which is ok to ignore - [Synth 8-2507] parameter declaration becomes local in MCycle with formal parameter declaration list...

    parameter COMPUTING = 1'b1 ; // this line will also cause the above warning
    reg state = IDLE ;
    reg n_state = IDLE ;
   
    reg done ;
    reg [7:0] count = 0 ; // assuming no computation takes more than 256 cycles.
    reg [2*width-1:0] temp_sum = 0 ;
    reg [2*width-1:0] shifted_op1 = 0 ;
    reg [2*width-1:0] shifted_op2 = 0 ;     
   
   //ADDED - For Both MCycle & Improved MCycle//
   reg Div_signed = 0;
   reg Neg_Op1 = 0;
   reg Neg_Op2 = 0;
   
  //ADDED - Improved MCycle -> Combinational Logic (Increase Hardware) to Cut cycles by up to n/2 cycles//
  //operand1_1, operand1_2 -> Multiplicant Left bit shift by 1 bit and by 2 bits 
  wire [2*width-1 : 0] operand1_1 = { shifted_op1[2*width-2 : 0], 1'b0 };       
  wire [2*width-1 : 0] operand1_2 = { shifted_op1[2*width-3 : 0], 2'b00 };      
  //operand2_1, operand2_2 -> Multiplier Right bit shift by 1 and by 2 bits
  wire [2*width-1 : 0] operand2_1 = { 1'b0, shifted_op2[2*width-1 : 1] };       
  wire [2*width-1 : 0] operand2_2 = { 2'b00, shifted_op2[2*width-1 : 2] };     
  //Determinine if LSB of Multiplier Op2 is 1 or 0 -> if 1 = Op1 taken as is, if 0, Check 2nd LSB if 1 or 0, if 1 take bit shifted Op1
  wire [2*width-1 : 0] next_value = shifted_op2[0] ? shifted_op1 : shifted_op2[1] ? operand1_1 : 0;
 //Compute new Sum
  wire [2*width-1 : 0] update_sum = temp_sum + next_value;
  //Update Op1 and Op2 based on the already shifted value of Op1 and Op2
  //next_operand is op1 bit shifted by 1 if op2 LSB was 1, if op2 is 0 return op1, 
  //else it would have mean 2nd LSB was 1 and next op1 is bit shifted twice
  //Similar logic for Op2
  wire [2*width-1 : 0] next_operand1 = shifted_op2[0] ? operand1_1 : 
                                       shifted_op2 == 0? shifted_op1 :
                                       operand1_2;
  wire [2*width-1 : 0] next_operand2 = shifted_op2[0] ? operand2_1 : 
                                       shifted_op2 == 0? shifted_op2 :
                                       operand2_2;
  
    always@( state, done, Start, RESET ) begin : IDLE_PROCESS  
		// Note : This block uses non-blocking assignments to get around an unpredictable Verilog simulation behaviour.
        // default outputs
        Busy <= 1'b0 ;
        n_state <= IDLE ;
        
        // reset
        if(~RESET)
            case(state)
                IDLE: begin
                    if(Start) begin // note: a mealy machine, since output depends on current state (IDLE) & input (Start)
                        n_state <= COMPUTING ;
                        Busy <= 1'b1 ;
                    end
                end
                COMPUTING: begin
                    if(~done) begin
                        n_state <= COMPUTING ;
                        Busy <= 1'b1 ;
                    end
                end        
            endcase    
    end


    always@( posedge CLK ) begin : STATE_UPDATE_PROCESS // state updating
        state <= n_state ;    
    end

    
    always@( posedge CLK ) begin : COMPUTING_PROCESS // process which does the actual computation
        // n_state == COMPUTING and state == IDLE implies we are just transitioning into COMPUTING
        done <= 1'b0 ; 
        if( RESET | (n_state == COMPUTING & state == IDLE) ) begin // 2nd condition is true during the very 1st clock cycle of the multiplication
            count = 0 ;
            temp_sum = 0 ;
            
            //MCycleOp - '00' Sign Mul, '01' Unsign Mul, '10' Sign Div, '11' Unsign Div
            //Check for Unsigned Division
            if (MCycleOp == 2'b11) begin
                shifted_op1 = { {width{1'b0}}, Operand1 };          //Dividend 0000...Dividend bits
                shifted_op2 = { Operand2, {width{1'b0}} };          //Divisor Divisor bits...0000
            end
            
            else begin
            shifted_op1 = { {width{~MCycleOp[0] & Operand1[width-1]}}, Operand1 } ; // sign extend the operand
            shifted_op2 = { {width{~MCycleOp[0] & Operand2[width-1]}}, Operand2 } ; 
            end
        end 
        
        //Pre Processing---------------------------------------------------------------------------------------------------------------------
        //Slide 24 - Conversion of Negative Operands to Positives before division -> Negate Result if Orignal Operands Different signs
        else if ( ~MCycleOp[0] & !Div_signed ) begin                       //Check if Sign Division Selected -> Serves as intermediate step for Sign Div
            //FOR MULTIPLICATION
            if (MCycleOp[1] == 0) begin
                if (shifted_op1[width-1] == 1) begin 
                    Neg_Op1 = 1;
                    shifted_op1 = ~(shifted_op1 - 1);                              //Converting NEG to POS Op1 - 2's Complement by -1 from original, Flip Op1             
                    Div_signed = 1;
                end
                if (shifted_op2[width-1] == 1) begin 
                    Neg_Op2 = 1;
                    shifted_op2 = ~(shifted_op2 - 1);                              //Converting NEG to POS Op2 - 2's Complement by -1 from original, Flip Op2                 
                    Div_signed = 1;
                end
            end    
            //FOR DIVISION
            else begin
                if (shifted_op1[width-1] == 1) begin                           //Op1 Dividend
                    Neg_Op1 = 1;
                    shifted_op1 = shifted_op1 - 1;                              //Converting NEG to POS Op1 - 2's Complement by -1 from original  (will flip in next step)
                    shifted_op1 = { {width{1'b0}}, ~shifted_op1[width-1:0] };   //Flip Op1 (2's Complement), 0000...Dividend bits                      
                    Div_signed = 1;
                end
                if (shifted_op2[width-1] == 1) begin                           //Op2 Divisor NEG
                    Neg_Op2 = 1;
                    shifted_op2 = shifted_op2 - 1;                             //Converting NEG to POS Op2 - 2's Complement by -1 from original (will flip in next step)
                    shifted_op2 = { ~shifted_op2[width-1:0], {width{1'b0}} };  //Flip Op2 (2's Complement), Divisor bits...0000
                    Div_signed = 1;
                end
                else begin 
                    shifted_op2 = { Operand2, {width{1'b0}} };                 //Op2 Divisor POS Divisor bits...0000
                end      
            end        
        end
        
        //Multiply---------------------------------------------------------------------------------------------------------------------
        //THIS WAS THE ORIGINAL GIVEN MULTIPLIER//
        //Sequential Multiplier - Slide 19
//        else if( ~MCycleOp[1] ) begin // Multiply
//            // if( ~MCycleOp[0] ), takes 2*'width' cycles to execute, returns signed(Operand1)*signed(Operand2)
//            // if( MCycleOp[0] ), takes 'width' cycles to execute, returns unsigned(Operand1)*unsigned(Operand2)        
            
//            //shifted_op2[0] is the multiplier Every cycle we check LSB of the Multiplier if 1, we add shifted Multiplicand
//            if( shifted_op2[0] ) // add only if b0 = 1
//                temp_sum = temp_sum + shifted_op1 ; // partial product for multiplication
            
//            //Here we bit right bit shift Op2 by 1 (Added 0 to MSB), left bit shift Op1 (Added 0 to LSB)
//            shifted_op2 = {1'b0, shifted_op2[2*width-1 : 1]} ;
//            shifted_op1 = {shifted_op1[2*width-2 : 0], 1'b0} ;    
            
//            //Track if Multiplication Completed
//            if( (MCycleOp[0] & count == width-1) | (~MCycleOp[0] & count == 2*width-1) ) // last cycle?
//                done <= 1'b1 ;   
               
//            count = count + 1;    
//        end    
          
          //NEW MULTIPLIER USING COMBINATIONAL LOGIC TO CONSIDER 2 LSB WORTH OF MULTIPLIER
        else if( ~MCycleOp[1] ) begin // Multiply
            //Update Values from Combinational Circuit
            shifted_op1 <= next_operand1;
            shifted_op2 <= next_operand2;
            temp_sum <= update_sum;
            //Once op1 and op2 (multiplicand and multiplier) are 0, done is set to 1
            done <= !(next_operand1 && next_operand2);
            //when not done -> flags are not cleared, once done -> flags cleared
            if (!done) begin
                Div_signed <= Div_signed;
                Neg_Op1 <= Neg_Op1;
                Neg_Op2 <= Neg_Op2;
            end
            else begin
                Div_signed <= 0;
                Neg_Op1 <= 0;
                Neg_Op2 <= 0;
            end
        end
        
        //Division--------------------------------------------------------------------------------------------------------------
        else if (MCycleOp[0] | Div_signed) begin
            //When Dividend < Divisor -> Quotient is 0, Remainder(Dividend) does not change till Division is carried out
            if (shifted_op1 < shifted_op2) begin                          
                //Remainder
                temp_sum[2*width-1 : width] = shifted_op1[width-1 : 0];    
                //Quotient - Shift left logic 0
                temp_sum[width-1 : 0] = {temp_sum[width-2 : 0], 1'b0};     
            end
            else begin                                                    
                //Once shifted_op2 aka Divisor Becomes Smaller or equal, do real division take place and Quotient =1  and Remainder changes
                shifted_op1 = shifted_op1 - shifted_op2;                  //Remainder - Divisor
                temp_sum[2*width-1: width] = shifted_op1[width-1 : 0];    //Store the above result into temp, Represent new 'Remainder' aka dividend
                temp_sum[width-1 : 0] = {temp_sum[width-2 : 0], 1'b1};    //Quotient Shift left logic 1
            end
            
            if (count == width) begin       //Flags reset at end of cycle
                done <= 1'b1;
                Neg_Op1 <= 0;
                Neg_Op2 <= 0;
                Div_signed <= 0;
            end
            else begin
                count = count + 1;
                shifted_op2 = { 1'b0, shifted_op2[2*width-1 : 1] };     //Divisor Shift Right
            end
        end
    end
    always @ (*) begin
                //Results--------------------------------------------------------------------------------------------------------------
            //Logic here is: Negate result if Operands were of Different Signs
            if (Neg_Op1 != Neg_Op2) begin
                Result2 = ~temp_sum[2*width-1 : width] + 1;
                Result1 = ~temp_sum[width-1 : 0] + 1 ;
            end
            else begin
                Result2 = temp_sum[2*width-1 : width] ;
                Result1 = temp_sum[width-1 : 0] ;
            end   
    end
endmodule

















