
----------------------------------------------------------------
-- Instruction Memory
----------------------------------------------------------------
constant INSTR_MEM : MEM_128x32 := (		x"E59F11F8", 
											x"E59F21F8", 
											x"E59F3214", 
											x"E5924000", 
											x"E5814000", 
											x"E2533001", 
											x"1AFFFFFD", 
											x"E1A0100F", 
											x"E59F0204", 
											x"E58F57D4", 
											x"E59F57D0", 
											x"E59F21F4", 
											x"E5820000", 
											x"E5820004", 
											x"EAFFFFFE", 
											others => x"00000000");

----------------------------------------------------------------
-- Data (Constant) Memory
----------------------------------------------------------------
constant DATA_CONST_MEM : MEM_128x32 := (	x"00000C00", 
											x"00000C04", 
											x"00000C08", 
											x"00000C0C", 
											x"00000C10", 
											x"00000C14", 
											x"00000C18", 
											x"00000000", 
											x"000000FF", 
											x"00000002", 
											x"00000800", 
											x"ABCD1234", 
											x"65570A0D", 
											x"6D6F636C", 
											x"6F742065", 
											x"33474320", 
											x"2E373032", 
											x"000A0D2E", 
											x"00000230", 
											others => x"00000000");

